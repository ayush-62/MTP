module test_obf ( line1, line2, reset, clock, outp, overflw );
  input line1, line2, reset, clock;
  output outp, overflw;
  wire   ____1, ____2, _____, _____0, ____, _______, _44, _42____, ___234,
         _43____, _41____, ___237, _108, _109, _110, _111, _112, _113, _114,
         _115, _116, _117, _118, _73, _323, _324, _325, _326, _327, _328, _329,
         _330, _331, _332, _333, _334, _335, _336, _337, _338, _339, _340,
         _341, _342, _343, _344, _345, _346, _347, _348, _349, _350, _351,
         _352, _353, _354, _355, _356, _357, _358, _359, _360, _361, _362,
         _363, _364, _365, _366, _367, _368, _369, _370, _371, _372, _373,
         _374, _375, _376, _377, _378, _379, _380, _381, _382, _383, _384,
         _385, _386, _387, _388, _389, _390, _391, _392, _393, _394, _395,
         _396, _397, _398, _399, _400, _401, _402, _403, _404, _405, _406,
         _407, _408, _409, _410, _411, _412, _413, _414, _415, _416, _417,
         _418, _419, _420, _421, _422, _423, _424, _425, _426, _427, _428,
         _429, _430, _431, _432, _433, _434, _435, _436, _437, _438, _439,
         _440, _441, _442, _443, _444, _445, _446, _447, _448, _449, _450,
         _451, _452, _453, _454, _455, _456, _457, _458, _459, _460, _461,
         _462, _463, _464, _465, _466, _467, _468, _469, _470, _471, _472,
         _473, _474, _475, _476, _477, _478, _479, _480, _481, _482, _483,
         _484, _485, _486, _487, _488, _489, _490, _491, _492, _493, _494,
         _495, _496, _497, _498, _499, _500, _501, _502, _503, _504, _505,
         _506, _507, _508, _509, _510, _511, _512, _513, _514, _515, _516,
         _517, _518, _519, _520, _521, _522, _523, _524, _525, _526, _527,
         _528, _529, _530, _531, _532, _533, _534, _535, _536, _537, _538,
         _539, _540, _541, _542, _543, _544, _545, _546, _547, _548, _549,
         _550, _551, _552, _553, _554, _555, _556, _557, _558, _559, _560,
         _561, _562, _563, _564, _565, _566, _567, _568, _569, _570, _571,
         _572, _573, _574, _575, _576, _577, _578, _579, _580, _581, _582,
         _583, _584, _585, _586, _587, _588, _589, _590, _591, _592, _593,
         _594, _595, _596, _597, _598, _599, _600, _601, _602, _603, _604,
         _605, _606, _607, _608, _609, _610, _611, _612, _613, _614, _615,
         _616, _617, _618, _619, _620, _621, _622, _623, _624, _625, _626,
         _627, _628, _629, _630, _631, _632, _633, _634, _635, _636, _637;
  wire   [10:0] ____0___________;
  assign ____1 = line1;
  assign ____2 = line2;
  assign _____ = reset;
  assign _____0 = clock;
  assign outp = ____;
  assign overflw = _______;

  dfrbp_1 ___________ ( .D(_323), .CLK(_____0), .RESET_B(_73), .Q(_______) );
  dfrbp_1 ________ ( .D(_44), .CLK(_____0), .RESET_B(_73), .Q(____) );
  dfxbp_1 ___________1_ ( .D(_42____), .CLK(_____0), .Q(_325), .Q_N(___234) );
  dfxbp_1 ___________2_ ( .D(_43____), .CLK(_____0), .Q(_324) );
  dfxbp_1 ___________0_ ( .D(_41____), .CLK(_____0), .Q_N(___237) );
  dfxtp_1 ____0________________0_ ( .D(_108), .CLK(_____0), .Q(
        ____0___________[0]) );
  dfxtp_1 ____0________________1_ ( .D(_109), .CLK(_____0), .Q(
        ____0___________[1]) );
  dfxtp_1 ____0________________5_ ( .D(_113), .CLK(_____0), .Q(
        ____0___________[5]) );
  dfxtp_1 ____0________________4_ ( .D(_112), .CLK(_____0), .Q(
        ____0___________[4]) );
  dfxtp_1 ____0________________3_ ( .D(_111), .CLK(_____0), .Q(
        ____0___________[3]) );
  dfxtp_1 ____0________________2_ ( .D(_110), .CLK(_____0), .Q(
        ____0___________[2]) );
  dfxtp_1 ____0________________10_ ( .D(_118), .CLK(_____0), .Q(
        ____0___________[10]) );
  dfxtp_1 ____0________________6_ ( .D(_114), .CLK(_____0), .Q(
        ____0___________[6]) );
  dfxtp_1 ____0________________7_ ( .D(_115), .CLK(_____0), .Q(
        ____0___________[7]) );
  dfxtp_1 ____0________________9_ ( .D(_117), .CLK(_____0), .Q(
        ____0___________[9]) );
  dfxtp_1 ____0________________8_ ( .D(_116), .CLK(_____0), .Q(
        ____0___________[8]) );
  xnor2_1 _341_inst ( .A(_326), .B(_327), .Y(_44) );
  nand2_1 _342_inst ( .A(_328), .B(_329), .Y(_327) );
  mux2i_1 _343_inst ( .A0(_330), .A1(_331), .S(_332), .Y(_43____) );
  nor2_1 _344_inst ( .A(_333), .B(_334), .Y(_332) );
  mux2i_1 _345_inst ( .A0(_335), .A1(_336), .S(_337), .Y(_334) );
  a21oi_1 _346_inst ( .A1(_338), .A2(_339), .B1(_____), .Y(_331) );
  o211ai_1 _347_inst ( .A1(_340), .A2(_328), .B1(_341), .C1(_342), .Y(_339) );
  o21ai_0 _348_inst ( .A1(_343), .A2(_344), .B1(_324), .Y(_338) );
  and2_0 _349_inst ( .A(____1), .B(_345), .X(_330) );
  o32ai_1 _350_inst ( .A1(_346), .A2(_347), .A3(_348), .B1(_349), .B2(_350), 
        .Y(_42____) );
  a21oi_1 _351_inst ( .A1(_347), .A2(_337), .B1(_345), .Y(_349) );
  a21oi_1 _352_inst ( .A1(___234), .A2(_351), .B1(_352), .Y(_348) );
  o32ai_1 _353_inst ( .A1(_353), .A2(_354), .A3(_355), .B1(_356), .B2(_357), 
        .Y(_352) );
  nor2_1 _354_inst ( .A(_343), .B(_324), .Y(_356) );
  o22ai_1 _355_inst ( .A1(_353), .A2(_328), .B1(_343), .B2(_355), .Y(_351) );
  inv_1 _356_inst ( .A(_329), .Y(_343) );
  inv_1 _357_inst ( .A(_335), .Y(_347) );
  nand2_1 _358_inst ( .A(____0___________[0]), .B(_336), .Y(_335) );
  mux2_1 _359_inst ( .A0(_358), .A1(_359), .S(_346), .X(_41____) );
  or3_1 _360_inst ( .A(_333), .B(_345), .C(_360), .X(_346) );
  inv_1 _361_inst ( .A(_361), .Y(_360) );
  o21ai_0 _362_inst ( .A1(____0___________[1]), .A2(_333), .B1(____1), .Y(_359) );
  a222oi_1 _363_inst ( .A1(_323), .A2(_329), .B1(_362), .B2(_73), .C1(_326), 
        .C2(_328), .Y(_358) );
  inv_1 _364_inst ( .A(_354), .Y(_328) );
  nor2_1 _365_inst ( .A(____1), .B(____2), .Y(_354) );
  nor2_1 _366_inst ( .A(_353), .B(_344), .Y(_326) );
  o32ai_1 _367_inst ( .A1(_363), .A2(_342), .A3(_325), .B1(_357), .B2(_329), 
        .Y(_362) );
  inv_1 _368_inst ( .A(_344), .Y(_357) );
  nor2_1 _369_inst ( .A(_341), .B(_340), .Y(_344) );
  xnor2_1 _370_inst ( .A(_340), .B(_329), .Y(_363) );
  inv_1 _371_inst ( .A(_355), .Y(_340) );
  nand2_1 _372_inst ( .A(____2), .B(____1), .Y(_329) );
  nor3_1 _373_inst ( .A(_355), .B(_342), .C(_341), .Y(_323) );
  a21oi_1 _374_inst ( .A1(_364), .A2(_365), .B1(_____), .Y(_118) );
  nor3_1 _375_inst ( .A(_366), .B(_367), .C(_368), .Y(_365) );
  o22ai_1 _376_inst ( .A1(_355), .A2(_369), .B1(_353), .B2(_370), .Y(_366) );
  nor3_1 _377_inst ( .A(_371), .B(_372), .C(_373), .Y(_364) );
  mux2i_1 _378_inst ( .A0(_374), .A1(_375), .S(_350), .Y(_371) );
  inv_1 _379_inst ( .A(_376), .Y(_375) );
  nor2_1 _380_inst ( .A(_377), .B(_378), .Y(_374) );
  a21oi_1 _381_inst ( .A1(_379), .A2(_380), .B1(_____), .Y(_117) );
  mux2i_1 _382_inst ( .A0(_381), .A1(_368), .S(_350), .Y(_380) );
  o21ai_0 _383_inst ( .A1(_353), .A2(_382), .B1(_383), .Y(_381) );
  nor2_1 _384_inst ( .A(_384), .B(_385), .Y(_379) );
  a21oi_1 _385_inst ( .A1(_386), .A2(_387), .B1(_____), .Y(_116) );
  mux2i_1 _386_inst ( .A0(_388), .A1(_389), .S(_350), .Y(_386) );
  or3_1 _387_inst ( .A(_390), .B(_377), .C(_391), .X(_389) );
  o32ai_1 _388_inst ( .A1(_392), .A2(_353), .A3(_393), .B1(_341), .B2(_394), 
        .Y(_391) );
  inv_1 _389_inst ( .A(_395), .Y(_393) );
  a21oi_1 _390_inst ( .A1(_396), .A2(_397), .B1(_____), .Y(_115) );
  nor3_1 _391_inst ( .A(_372), .B(_377), .C(_378), .Y(_397) );
  nand4_1 _392_inst ( .A(_398), .B(_399), .C(_400), .D(_401), .Y(_372) );
  nor3_1 _393_inst ( .A(_402), .B(_403), .C(_404), .Y(_401) );
  mux2i_1 _394_inst ( .A0(_405), .A1(_406), .S(_350), .Y(_402) );
  and3_1 _395_inst ( .A(_407), .B(_408), .C(_409), .X(_406) );
  nor2_1 _396_inst ( .A(_410), .B(_411), .Y(_405) );
  inv_1 _397_inst ( .A(_412), .Y(_398) );
  nor2_1 _398_inst ( .A(_376), .B(_413), .Y(_396) );
  mux2i_1 _399_inst ( .A0(_414), .A1(_415), .S(_350), .Y(_413) );
  and2_0 _400_inst ( .A(_416), .B(_383), .X(_415) );
  nor2_1 _401_inst ( .A(_367), .B(_417), .Y(_383) );
  inv_1 _402_inst ( .A(_368), .Y(_414) );
  nand3_1 _403_inst ( .A(_418), .B(_419), .C(_420), .Y(_368) );
  nand3_1 _404_inst ( .A(_421), .B(_422), .C(_423), .Y(_376) );
  a21oi_1 _405_inst ( .A1(_424), .A2(_425), .B1(_____), .Y(_114) );
  and4_1 _406_inst ( .A(_426), .B(_409), .C(_427), .D(_382), .X(_425) );
  nor2_1 _407_inst ( .A(_388), .B(_428), .Y(_426) );
  inv_1 _408_inst ( .A(_422), .Y(_388) );
  nor4_1 _409_inst ( .A(_377), .B(_429), .C(_384), .D(_430), .Y(_424) );
  mux2i_1 _410_inst ( .A0(_431), .A1(_432), .S(_350), .Y(_430) );
  nor4_1 _411_inst ( .A(_433), .B(_434), .C(_435), .D(_410), .Y(_432) );
  inv_1 _412_inst ( .A(_436), .Y(_435) );
  nand3_1 _413_inst ( .A(_437), .B(_438), .C(_439), .Y(_434) );
  nand4_1 _414_inst ( .A(_440), .B(_441), .C(_442), .D(_418), .Y(_433) );
  nor4_1 _415_inst ( .A(_443), .B(_444), .C(_445), .D(_446), .Y(_431) );
  inv_1 _416_inst ( .A(_447), .Y(_445) );
  o21ai_0 _417_inst ( .A1(_353), .A2(_448), .B1(_421), .Y(_444) );
  nand3_1 _418_inst ( .A(_408), .B(_449), .C(_450), .Y(_443) );
  and3_1 _419_inst ( .A(_451), .B(_369), .C(_452), .X(_450) );
  nand2_1 _420_inst ( .A(_453), .B(_454), .Y(_384) );
  mux2i_1 _421_inst ( .A0(_373), .A1(_390), .S(_350), .Y(_453) );
  inv_1 _422_inst ( .A(_455), .Y(_390) );
  a21oi_1 _423_inst ( .A1(_456), .A2(_457), .B1(_____), .Y(_113) );
  and4_1 _424_inst ( .A(_439), .B(_458), .C(_459), .D(_460), .X(_457) );
  nor3_1 _425_inst ( .A(_461), .B(_373), .C(_462), .Y(_456) );
  mux2i_1 _426_inst ( .A0(_463), .A1(_464), .S(_350), .Y(_461) );
  nor4_1 _427_inst ( .A(_465), .B(_466), .C(_467), .D(_468), .Y(_464) );
  nand3_1 _428_inst ( .A(_422), .B(_469), .C(_470), .Y(_466) );
  nand4_1 _429_inst ( .A(_471), .B(_472), .C(_418), .D(_473), .Y(_465) );
  and3_1 _430_inst ( .A(_474), .B(_475), .C(_370), .X(_473) );
  nor4_1 _431_inst ( .A(_476), .B(_477), .C(_478), .D(_479), .Y(_463) );
  nand3_1 _432_inst ( .A(_452), .B(_427), .C(_409), .Y(_477) );
  nand4_1 _433_inst ( .A(_480), .B(_440), .C(_481), .D(_482), .Y(_476) );
  and4_1 _434_inst ( .A(_483), .B(_484), .C(_420), .D(_485), .X(_440) );
  and3_1 _435_inst ( .A(_486), .B(_487), .C(_488), .X(_485) );
  and3_1 _436_inst ( .A(_489), .B(_490), .C(_491), .X(_420) );
  inv_1 _437_inst ( .A(_492), .Y(_480) );
  a21oi_1 _438_inst ( .A1(_493), .A2(_494), .B1(_____), .Y(_112) );
  and4_1 _439_inst ( .A(_495), .B(_370), .C(_496), .D(_497), .X(_494) );
  and2_0 _440_inst ( .A(_486), .B(_408), .X(_495) );
  nor4_1 _441_inst ( .A(_498), .B(_499), .C(_500), .D(_373), .Y(_493) );
  inv_1 _442_inst ( .A(_441), .Y(_500) );
  nand2_1 _443_inst ( .A(_501), .B(_502), .Y(_498) );
  inv_1 _444_inst ( .A(_503), .Y(_502) );
  mux2i_1 _445_inst ( .A0(_504), .A1(_492), .S(_350), .Y(_501) );
  nand2_1 _446_inst ( .A(_505), .B(_506), .Y(_492) );
  nand4_1 _447_inst ( .A(_487), .B(_427), .C(_394), .D(_507), .Y(_504) );
  inv_1 _448_inst ( .A(_508), .Y(_507) );
  o211ai_1 _449_inst ( .A1(_451), .A2(_355), .B1(_509), .C1(_474), .Y(_508) );
  nor2_1 _450_inst ( .A(_____), .B(_510), .Y(_111) );
  nor4_1 _451_inst ( .A(_511), .B(_512), .C(_499), .D(_513), .Y(_510) );
  mux2i_1 _452_inst ( .A0(_514), .A1(_515), .S(_350), .Y(_513) );
  nor4_1 _453_inst ( .A(_516), .B(_517), .C(_377), .D(_518), .Y(_515) );
  inv_1 _454_inst ( .A(_470), .Y(_377) );
  nand3_1 _455_inst ( .A(_451), .B(_496), .C(_486), .Y(_516) );
  nor4_1 _456_inst ( .A(_519), .B(_520), .C(_428), .D(_479), .Y(_514) );
  inv_1 _457_inst ( .A(_521), .Y(_479) );
  inv_1 _458_inst ( .A(_522), .Y(_428) );
  nand4_1 _459_inst ( .A(_409), .B(_436), .C(_370), .D(_475), .Y(_519) );
  nand4_1 _460_inst ( .A(_523), .B(_491), .C(_524), .D(_525), .Y(_499) );
  and3_1 _461_inst ( .A(_489), .B(_382), .C(_447), .X(_525) );
  mux2i_1 _462_inst ( .A0(_526), .A1(_527), .S(_350), .Y(_524) );
  nand4_1 _463_inst ( .A(_528), .B(_449), .C(_490), .D(_529), .Y(_527) );
  and4_1 _464_inst ( .A(_437), .B(_369), .C(_472), .D(_530), .X(_529) );
  nand4_1 _465_inst ( .A(_471), .B(_488), .C(_531), .D(_438), .Y(_526) );
  inv_1 _466_inst ( .A(_404), .Y(_523) );
  nand4_1 _467_inst ( .A(_532), .B(_439), .C(_455), .D(_452), .Y(_404) );
  o21ai_0 _468_inst ( .A1(_355), .A2(_496), .B1(_533), .Y(_512) );
  inv_1 _469_inst ( .A(_403), .Y(_533) );
  nand4_1 _470_inst ( .A(_418), .B(_505), .C(_422), .D(_534), .Y(_511) );
  nor2_1 _471_inst ( .A(_535), .B(_536), .Y(_534) );
  a21oi_1 _472_inst ( .A1(_537), .A2(_387), .B1(_____), .Y(_110) );
  and4_1 _473_inst ( .A(_538), .B(_539), .C(_454), .D(_540), .X(_387) );
  and4_1 _474_inst ( .A(_541), .B(_506), .C(_497), .D(_542), .X(_454) );
  nor2_1 _475_inst ( .A(_543), .B(_544), .Y(_542) );
  mux2i_1 _476_inst ( .A0(_505), .A1(_474), .S(_350), .Y(_544) );
  inv_1 _477_inst ( .A(_481), .Y(_543) );
  nand3_1 _478_inst ( .A(_545), .B(_546), .C(_547), .Y(_497) );
  inv_1 _479_inst ( .A(_385), .Y(_539) );
  nand3_1 _480_inst ( .A(_548), .B(_441), .C(_549), .Y(_385) );
  nor3_1 _481_inst ( .A(_536), .B(_520), .C(_467), .Y(_549) );
  inv_1 _482_inst ( .A(_483), .Y(_520) );
  inv_1 _483_inst ( .A(_459), .Y(_536) );
  nand3_1 _484_inst ( .A(_550), .B(_545), .C(_547), .Y(_441) );
  mux2_1 _485_inst ( .A0(_427), .A1(_530), .S(____1), .X(_548) );
  mux2i_1 _486_inst ( .A0(_551), .A1(_378), .S(_350), .Y(_538) );
  nand3_1 _487_inst ( .A(_482), .B(_442), .C(_484), .Y(_378) );
  nand2_1 _488_inst ( .A(_421), .B(_552), .Y(_551) );
  mux2i_1 _489_inst ( .A0(_553), .A1(_554), .S(_350), .Y(_537) );
  nand4_1 _490_inst ( .A(_419), .B(_458), .C(_490), .D(_555), .Y(_554) );
  a21oi_1 _491_inst ( .A1(_556), .A2(_557), .B1(_558), .Y(_555) );
  or3_1 _492_inst ( .A(_559), .B(_373), .C(_560), .X(_553) );
  o211ai_1 _493_inst ( .A1(_452), .A2(_353), .B1(_472), .C1(_469), .Y(_560) );
  inv_1 _494_inst ( .A(_342), .Y(_353) );
  nor2_1 _495_inst ( .A(_324), .B(_____), .Y(_342) );
  inv_1 _496_inst ( .A(_416), .Y(_373) );
  o21ai_0 _497_inst ( .A1(_487), .A2(_355), .B1(_407), .Y(_559) );
  a21oi_1 _498_inst ( .A1(_561), .A2(_562), .B1(_____), .Y(_109) );
  and4_1 _499_inst ( .A(_563), .B(_452), .C(_531), .D(_506), .X(_562) );
  nand3_1 _500_inst ( .A(_550), .B(_564), .C(_547), .Y(_506) );
  nor2_1 _501_inst ( .A(_518), .B(_558), .Y(_563) );
  inv_1 _502_inst ( .A(_489), .Y(_558) );
  inv_1 _503_inst ( .A(_442), .Y(_518) );
  nor4_1 _504_inst ( .A(_412), .B(_565), .C(_503), .D(_566), .Y(_561) );
  mux2i_1 _505_inst ( .A0(_567), .A1(_568), .S(_350), .Y(_566) );
  nor4_1 _506_inst ( .A(_446), .B(_569), .C(_367), .D(_517), .Y(_568) );
  nand3_1 _507_inst ( .A(_484), .B(_408), .C(_509), .Y(_517) );
  nor3_1 _508_inst ( .A(_478), .B(_410), .C(_467), .Y(_509) );
  and2_0 _509_inst ( .A(_570), .B(_336), .X(_467) );
  inv_1 _510_inst ( .A(_458), .Y(_410) );
  nand2_1 _511_inst ( .A(_469), .B(_522), .Y(_367) );
  nand2_1 _512_inst ( .A(_439), .B(_369), .Y(_569) );
  inv_1 _513_inst ( .A(_419), .Y(_446) );
  nor4_1 _514_inst ( .A(_571), .B(_572), .C(_573), .D(_556), .Y(_567) );
  inv_1 _515_inst ( .A(_532), .Y(_556) );
  inv_1 _516_inst ( .A(_491), .Y(_572) );
  nand2_1 _517_inst ( .A(_574), .B(_575), .Y(_491) );
  nand3_1 _518_inst ( .A(_459), .B(_482), .C(_400), .Y(_571) );
  and3_1 _519_inst ( .A(_451), .B(_475), .C(_488), .X(_400) );
  nand3_1 _520_inst ( .A(_546), .B(_564), .C(_547), .Y(_459) );
  and2_0 _521_inst ( .A(_576), .B(____0___________[6]), .X(_547) );
  nand2_1 _522_inst ( .A(_577), .B(_541), .Y(_503) );
  nand3_1 _523_inst ( .A(_546), .B(_564), .C(_578), .Y(_541) );
  mux2i_1 _524_inst ( .A0(_579), .A1(_580), .S(_350), .Y(_577) );
  inv_1 _525_inst ( .A(____1), .Y(_350) );
  nand4_1 _526_inst ( .A(_481), .B(_483), .C(_581), .D(_422), .Y(_580) );
  nand3_1 _527_inst ( .A(_550), .B(_564), .C(_578), .Y(_483) );
  nand2_1 _528_inst ( .A(_570), .B(____0___________[1]), .Y(_481) );
  and3_1 _529_inst ( .A(_545), .B(____0___________[3]), .C(_578), .X(_570) );
  and2_0 _530_inst ( .A(_576), .B(_582), .X(_578) );
  and4_1 _531_inst ( .A(____0___________[8]), .B(____0___________[2]), .C(
        ____0___________[9]), .D(_583), .X(_576) );
  nor3_1 _532_inst ( .A(____0___________[0]), .B(____0___________[7]), .C(
        ____0___________[10]), .Y(_583) );
  nand4_1 _533_inst ( .A(_540), .B(_418), .C(_399), .D(_448), .Y(_579) );
  o21ai_0 _534_inst ( .A1(_355), .A2(_475), .B1(_407), .Y(_565) );
  inv_1 _535_inst ( .A(_468), .Y(_407) );
  nand2_1 _536_inst ( .A(_447), .B(_528), .Y(_468) );
  nand2_1 _537_inst ( .A(___237), .B(_73), .Y(_355) );
  inv_1 _538_inst ( .A(_____), .Y(_73) );
  nand4_1 _539_inst ( .A(_438), .B(_487), .C(_530), .D(_584), .Y(_412) );
  inv_1 _540_inst ( .A(_585), .Y(_584) );
  o211ai_1 _541_inst ( .A1(_472), .A2(____1), .B1(_586), .C1(_471), .Y(_585)
         );
  nand3_1 _542_inst ( .A(_575), .B(_587), .C(_550), .Y(_487) );
  o21ai_0 _543_inst ( .A1(_588), .A2(_589), .B1(_395), .Y(_438) );
  a21oi_1 _544_inst ( .A1(_590), .A2(_591), .B1(_____), .Y(_108) );
  nor2_1 _545_inst ( .A(_592), .B(_593), .Y(_591) );
  nand4_1 _546_inst ( .A(_490), .B(_419), .C(_458), .D(_447), .Y(_593) );
  nand2_1 _547_inst ( .A(_594), .B(_595), .Y(_447) );
  nand3_1 _548_inst ( .A(_596), .B(_546), .C(_597), .Y(_458) );
  nand2_1 _549_inst ( .A(_598), .B(_599), .Y(_419) );
  nand3_1 _550_inst ( .A(_600), .B(_601), .C(_602), .Y(_490) );
  nand4_1 _551_inst ( .A(_530), .B(_472), .C(_452), .D(_475), .Y(_592) );
  nand2_1 _552_inst ( .A(_597), .B(_603), .Y(_475) );
  nand2_1 _553_inst ( .A(_575), .B(_604), .Y(_452) );
  nand3_1 _554_inst ( .A(_605), .B(_596), .C(_550), .Y(_472) );
  nand3_1 _555_inst ( .A(_602), .B(_600), .C(____0___________[5]), .Y(_530) );
  and4_1 _556_inst ( .A(_606), .B(_607), .C(_423), .D(_416), .X(_590) );
  a21oi_1 _557_inst ( .A1(_608), .A2(_595), .B1(_573), .Y(_416) );
  and3_1 _558_inst ( .A(_600), .B(_601), .C(_609), .X(_573) );
  and3_1 _559_inst ( .A(_370), .B(_369), .C(_552), .X(_423) );
  inv_1 _560_inst ( .A(_429), .Y(_552) );
  nand2_1 _561_inst ( .A(_521), .B(_531), .Y(_429) );
  nand3_1 _562_inst ( .A(____0___________[5]), .B(_609), .C(_610), .Y(_531) );
  nand3_1 _563_inst ( .A(_611), .B(_546), .C(_612), .Y(_521) );
  nand2_1 _564_inst ( .A(_589), .B(_597), .Y(_369) );
  nand2_1 _565_inst ( .A(_613), .B(_614), .Y(_370) );
  mux2_1 _566_inst ( .A0(_615), .A1(_616), .S(____1), .X(_607) );
  nor4_1 _567_inst ( .A(_617), .B(_618), .C(_411), .D(_619), .Y(_616) );
  inv_1 _568_inst ( .A(_418), .Y(_619) );
  nand4_1 _569_inst ( .A(_597), .B(_550), .C(_602), .D(_620), .Y(_418) );
  inv_1 _570_inst ( .A(_486), .Y(_411) );
  nand3_1 _571_inst ( .A(_550), .B(_596), .C(_597), .Y(_486) );
  nand3_1 _572_inst ( .A(_439), .B(_455), .C(_528), .Y(_618) );
  nand2_1 _573_inst ( .A(_599), .B(_621), .Y(_528) );
  nand3_1 _574_inst ( .A(_596), .B(_546), .C(_605), .Y(_455) );
  and2_0 _575_inst ( .A(_611), .B(_602), .X(_596) );
  nand2_1 _576_inst ( .A(_395), .B(_604), .Y(_439) );
  nand4_1 _577_inst ( .A(_421), .B(_586), .C(_470), .D(_469), .Y(_617) );
  nand3_1 _578_inst ( .A(_620), .B(____0___________[1]), .C(_598), .Y(_469) );
  nand2_1 _579_inst ( .A(_599), .B(_595), .Y(_470) );
  and2_0 _580_inst ( .A(_611), .B(____0___________[1]), .X(_599) );
  and4_1 _581_inst ( .A(_460), .B(_505), .C(_436), .D(_449), .X(_586) );
  nand2_1 _582_inst ( .A(_614), .B(_603), .Y(_449) );
  nand2_1 _583_inst ( .A(_589), .B(_605), .Y(_436) );
  nand4_1 _584_inst ( .A(_605), .B(_546), .C(_609), .D(_620), .Y(_505) );
  and4_1 _585_inst ( .A(_382), .B(_394), .C(_437), .D(_496), .X(_460) );
  nand2_1 _586_inst ( .A(_603), .B(_395), .Y(_496) );
  nand2_1 _587_inst ( .A(_613), .B(_395), .Y(_394) );
  nand2_1 _588_inst ( .A(_613), .B(_597), .Y(_382) );
  nor2_1 _589_inst ( .A(_535), .B(_478), .Y(_421) );
  and2_0 _590_inst ( .A(_621), .B(_608), .X(_478) );
  inv_1 _591_inst ( .A(_581), .Y(_535) );
  nand2_1 _592_inst ( .A(_598), .B(_608), .Y(_581) );
  and2_0 _593_inst ( .A(_622), .B(_564), .X(_598) );
  nor4_1 _594_inst ( .A(_623), .B(_624), .C(_417), .D(_462), .Y(_615) );
  nand4_1 _595_inst ( .A(_442), .B(_408), .C(_532), .D(_399), .Y(_462) );
  nand3_1 _596_inst ( .A(_604), .B(_582), .C(_545), .Y(_399) );
  and2_0 _597_inst ( .A(_546), .B(_587), .X(_604) );
  nand2_1 _598_inst ( .A(_588), .B(_575), .Y(_532) );
  nor3_1 _599_inst ( .A(____0___________[4]), .B(____0___________[5]), .C(_582), .Y(_575) );
  inv_1 _600_inst ( .A(_392), .Y(_588) );
  nand3_1 _601_inst ( .A(____0___________[5]), .B(_602), .C(_610), .Y(_408) );
  nand2_1 _602_inst ( .A(_621), .B(_594), .Y(_442) );
  and2_0 _603_inst ( .A(_622), .B(_545), .X(_621) );
  inv_1 _604_inst ( .A(_540), .Y(_417) );
  nand3_1 _605_inst ( .A(_546), .B(_620), .C(_612), .Y(_540) );
  nor2_1 _606_inst ( .A(____0___________[1]), .B(____0___________[3]), .Y(_546) );
  nand3_1 _607_inst ( .A(_422), .B(_522), .C(_482), .Y(_624) );
  nand4_1 _608_inst ( .A(_605), .B(_608), .C(_609), .D(_625), .Y(_482) );
  nand3_1 _609_inst ( .A(_545), .B(____0___________[6]), .C(_574), .Y(_522) );
  and3_1 _610_inst ( .A(_602), .B(____0___________[3]), .C(_608), .X(_574) );
  nand3_1 _611_inst ( .A(_608), .B(_625), .C(_612), .Y(_422) );
  and3_1 _612_inst ( .A(_626), .B(_627), .C(_333), .X(_608) );
  nand4_1 _613_inst ( .A(_489), .B(_409), .C(_628), .D(_471), .Y(_623) );
  nand3_1 _614_inst ( .A(_629), .B(_582), .C(_545), .Y(_471) );
  nor2_1 _615_inst ( .A(_601), .B(____0___________[4]), .Y(_545) );
  o21ai_0 _616_inst ( .A1(_630), .A2(_631), .B1(_392), .Y(_629) );
  nand2_1 _617_inst ( .A(_632), .B(_625), .Y(_392) );
  inv_1 _618_inst ( .A(_550), .Y(_631) );
  and2_0 _619_inst ( .A(_451), .B(_488), .X(_628) );
  nand2_1 _620_inst ( .A(_589), .B(_614), .Y(_488) );
  and2_0 _621_inst ( .A(_564), .B(_582), .X(_614) );
  nand2_1 _622_inst ( .A(_603), .B(_605), .Y(_451) );
  and2_0 _623_inst ( .A(_632), .B(____0___________[3]), .X(_603) );
  and2_0 _624_inst ( .A(_633), .B(_345), .X(_632) );
  nor3_1 _625_inst ( .A(____0___________[0]), .B(____0___________[2]), .C(_336), .Y(_345) );
  nand3_1 _626_inst ( .A(_550), .B(_611), .C(_612), .Y(_409) );
  and2_0 _627_inst ( .A(_597), .B(_609), .X(_612) );
  nor3_1 _628_inst ( .A(____0___________[5]), .B(____0___________[6]), .C(
        ____0___________[4]), .Y(_597) );
  nand3_1 _629_inst ( .A(_609), .B(_601), .C(_610), .Y(_489) );
  and4_1 _630_inst ( .A(_620), .B(_634), .C(____0___________[1]), .D(_635), 
        .X(_610) );
  a211oi_1 _631_inst ( .A1(_395), .A2(_589), .B1(_403), .C1(_636), .Y(_606) );
  o21ai_0 _632_inst ( .A1(_437), .A2(_341), .B1(_484), .Y(_636) );
  nand3_1 _633_inst ( .A(_609), .B(_600), .C(____0___________[5]), .Y(_484) );
  and4_1 _634_inst ( .A(_620), .B(_634), .C(_336), .D(_635), .X(_600) );
  nor3_1 _635_inst ( .A(_626), .B(_361), .C(_627), .Y(_620) );
  inv_1 _636_inst ( .A(____0___________[8]), .Y(_627) );
  inv_1 _637_inst ( .A(_557), .Y(_341) );
  nor2_1 _638 ( .A(_____), .B(___234), .Y(_557) );
  nand2_1 _639 ( .A(_613), .B(_605), .Y(_437) );
  nor3_1 _640 ( .A(_635), .B(_582), .C(_601), .Y(_605) );
  nor3_1 _641 ( .A(_625), .B(____0___________[1]), .C(_630), .Y(_613) );
  nand3_1 _642 ( .A(_448), .B(_427), .C(_474), .Y(_403) );
  nand3_1 _643 ( .A(_595), .B(_336), .C(_611), .Y(_474) );
  nor3_1 _644 ( .A(____0___________[7]), .B(____0___________[8]), .C(_361), 
        .Y(_611) );
  nand2_1 _645 ( .A(____0___________[2]), .B(____0___________[0]), .Y(_361) );
  and3_1 _646 ( .A(_564), .B(_634), .C(_602), .X(_595) );
  and2_0 _647 ( .A(____0___________[9]), .B(____0___________[10]), .X(_602) );
  nor2_1 _648 ( .A(_635), .B(____0___________[5]), .Y(_564) );
  nand4_1 _649 ( .A(_622), .B(_594), .C(_635), .D(_601), .Y(_427) );
  and3_1 _650 ( .A(____0___________[8]), .B(____0___________[7]), .C(_333), 
        .X(_594) );
  nor3_1 _651 ( .A(____0___________[1]), .B(____0___________[2]), .C(
        ____0___________[0]), .Y(_333) );
  and2_0 _652 ( .A(_609), .B(_634), .X(_622) );
  nor2_1 _653 ( .A(_582), .B(_625), .Y(_634) );
  inv_1 _654 ( .A(____0___________[6]), .Y(_582) );
  nor2_1 _655 ( .A(____0___________[10]), .B(____0___________[9]), .Y(_609) );
  nand3_1 _656 ( .A(_395), .B(_587), .C(_550), .Y(_448) );
  nor2_1 _657 ( .A(_336), .B(____0___________[3]), .Y(_550) );
  inv_1 _658 ( .A(_630), .Y(_587) );
  nor3_1 _659 ( .A(_625), .B(_336), .C(_630), .Y(_589) );
  nand3_1 _660 ( .A(____0___________[0]), .B(_337), .C(_633), .Y(_630) );
  nor4_1 _661 ( .A(_637), .B(_626), .C(____0___________[8]), .D(
        ____0___________[9]), .Y(_633) );
  inv_1 _662 ( .A(____0___________[7]), .Y(_626) );
  inv_1 _663 ( .A(____0___________[10]), .Y(_637) );
  inv_1 _664 ( .A(____0___________[2]), .Y(_337) );
  inv_1 _665 ( .A(____0___________[1]), .Y(_336) );
  inv_1 _666 ( .A(____0___________[3]), .Y(_625) );
  nor3_1 _667 ( .A(_635), .B(____0___________[6]), .C(_601), .Y(_395) );
  inv_1 _668 ( .A(____0___________[5]), .Y(_601) );
  inv_1 _669 ( .A(____0___________[4]), .Y(_635) );
endmodule

