module test_org ( line1, line2, reset, outp, overflw, clock );
  input line1, line2, reset, clock;
  output outp, overflw;
  wire   N41, N42, n1, n2, n3, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50;
  wire   [2:0] stato;

  dfrtp_1 \stato_reg[0]  ( .D(N41), .CLK(clock), .RESET_B(n1), .Q(stato[0]) );
  dfrtp_1 \stato_reg[1]  ( .D(N42), .CLK(clock), .RESET_B(n1), .Q(stato[1]) );
  dfrtp_1 \stato_reg[2]  ( .D(n2), .CLK(clock), .RESET_B(n1), .Q(stato[2]) );
  dfrtp_1 overflw_reg ( .D(n3), .CLK(clock), .RESET_B(n1), .Q(overflw) );
  dfrtp_1 outp_reg ( .D(n28), .CLK(clock), .RESET_B(n1), .Q(outp) );
  xor2_1 U33 ( .A(n29), .B(n30), .X(n28) );
  nand2_1 U34 ( .A(stato[2]), .B(n31), .Y(n30) );
  o22ai_1 U35 ( .A1(stato[2]), .A2(n32), .B1(stato[1]), .B2(n33), .Y(n2) );
  nor2_1 U36 ( .A(n34), .B(n35), .Y(n33) );
  a21oi_1 U37 ( .A1(n36), .A2(n29), .B1(n37), .Y(n34) );
  nor2_1 U38 ( .A(n38), .B(n35), .Y(n32) );
  inv_1 U39 ( .A(reset), .Y(n1) );
  o221ai_1 U40 ( .A1(n36), .A2(n39), .B1(n40), .B2(n37), .C1(n41), .Y(N42) );
  o21ai_0 U41 ( .A1(n35), .A2(n37), .B1(n38), .Y(n41) );
  a21oi_1 U42 ( .A1(n42), .A2(n29), .B1(n43), .Y(n40) );
  a21oi_1 U43 ( .A1(n44), .A2(n29), .B1(n36), .Y(n43) );
  nand2_1 U44 ( .A(n45), .B(n46), .Y(N41) );
  mux2i_1 U45 ( .A0(n47), .A1(n48), .S(n37), .Y(n46) );
  nor2_1 U46 ( .A(stato[0]), .B(n39), .Y(n48) );
  inv_1 U47 ( .A(n42), .Y(n39) );
  nor2_1 U48 ( .A(n35), .B(stato[1]), .Y(n42) );
  inv_1 U49 ( .A(n44), .Y(n35) );
  nor2_1 U50 ( .A(n38), .B(n29), .Y(n47) );
  o21ai_0 U51 ( .A1(line2), .A2(line1), .B1(n44), .Y(n29) );
  mux2i_1 U52 ( .A0(n49), .A1(n3), .S(n44), .Y(n45) );
  nand2_1 U53 ( .A(line2), .B(line1), .Y(n44) );
  nor3_1 U54 ( .A(n36), .B(stato[2]), .C(n50), .Y(n3) );
  o211ai_1 U55 ( .A1(stato[1]), .A2(n36), .B1(n31), .C1(n37), .Y(n49) );
  inv_1 U56 ( .A(stato[2]), .Y(n37) );
  inv_1 U57 ( .A(n38), .Y(n31) );
  nor2_1 U58 ( .A(n50), .B(stato[0]), .Y(n38) );
  inv_1 U59 ( .A(stato[1]), .Y(n50) );
  inv_1 U60 ( .A(stato[0]), .Y(n36) );
endmodule

