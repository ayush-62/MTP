`timescale 1ns / 1ps


module toy_obf ( datain, clk, rst, op, valid, dataout );
  input [7:0] datain;
  input [1:0] op;
  output [7:0] dataout;
  input clk, rst;
  output valid;
  wire   ___0____1999, ___0____1998, ___0____2003, ___0_0__1996, ___0____1997,
         ___0____2004, ___0____1994, ___0_9__1995, ___09___2017, ___0____1991,
         ___0____1992, ___0____2008, ___0____2007, ___0____1990, ___0____2005,
         ___0____1987, ___0____1989, ___0____2006, ___0____1983, ___0____1985,
         ___0____1982, ___0____1981, __99___1933, __99___1932, __9____1926,
         __9____1920, __9____1899, __9____1911, __9____1887, __9____1882,
         __9_9__1884, __9____1881, __9____1869, __9____1860, __9_9,
         __9____1861, __9____1872, __9____1870, __9____1868, __9____1873,
         __90___1854, __90_, ___99__1850, ____0___2025, _______________1154,
         _______1827, _______1830, _______1826, ___09___2013, _______1828,
         _______1820, ____0__1814, _______1806, _______1801, _______1793,
         _______1798, _______1794, _______1781, ___________0___1152,
         ___0___1764, _______1652, _______1397, n2, n45, n47, n48, n124, n125,
         n159, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033;

  dfxbp_1 _______________ ( .D(___0____1999), .CLK(clk), .Q(dataout[5]) );
  dfxbp_1 _______________36111 ( .D(___0____1998), .CLK(clk), .Q(dataout[4])
         );
  dfxbp_1 _______________36112 ( .D(___0_0__1996), .CLK(clk), .Q(dataout[1])
         );
  dfxbp_1 _____________0_ ( .D(___0____1997), .CLK(clk), .Q(dataout[0]) );
  dfxbp_1 _______________36113 ( .D(___0____1994), .CLK(clk), .Q_N(dataout[7])
         );
  dfxbp_1 _______________36114 ( .D(___0_9__1995), .CLK(clk), .Q_N(dataout[6])
         );
  dfxbp_1 ____________ ( .D(___09___2017), .CLK(clk), .Q_N(___0____2003) );
  dfxbp_1 _______________36115 ( .D(___0____1991), .CLK(clk), .Q(dataout[2])
         );
  dfxbp_1 _______________36116 ( .D(___0____1992), .CLK(clk), .Q(dataout[3])
         );
  dfxbp_1 ____________36117 ( .D(___0____1990), .CLK(clk), .Q_N(___0____2004)
         );
  dfxbp_1 ____________36118 ( .D(___0____1987), .CLK(clk), .Q_N(___0____2007)
         );
  dfxbp_1 __________0_ ( .D(___0____1989), .CLK(clk), .Q_N(___0____2008) );
  dfxbp_1 ____________36120 ( .D(___0____1983), .CLK(clk), .Q(n124) );
  dfxbp_1 ____________36121 ( .D(___0____1985), .CLK(clk), .Q(n125) );
  dfxbp_1 ____________36122 ( .D(___0____1982), .CLK(clk), .Q_N(___0____2006)
         );
  dfxbp_1 ____________36123 ( .D(___0____1981), .CLK(clk), .Q_N(___0____2005)
         );
  dfxbp_1 __________________ ( .D(__99___1933), .CLK(clk), .Q(n1016), .Q_N(
        n538) );
  dfxbp_1 ________0_ ( .D(__99___1932), .CLK(clk), .Q(n1014) );
  dfrbp_1 __________________36151 ( .D(n45), .CLK(clk), .RESET_B(rst), .Q_N(
        n1023) );
  dfxbp_1 __________________36155 ( .D(__9____1926), .CLK(clk), .Q(n1027), 
        .Q_N(n539) );
  dfrbp_1 __________________36160 ( .D(__9____1920), .CLK(clk), .RESET_B(rst), 
        .Q(n532), .Q_N(n1020) );
  dfrbp_1 _______________________ ( .D(__9____1899), .CLK(clk), .RESET_B(rst), 
        .Q(n997), .Q_N(n522) );
  dfrbp_1 _______________________36161 ( .D(__9____1911), .CLK(clk), .RESET_B(
        rst), .Q(n998), .Q_N(n517) );
  dfxbp_1 __________ ( .D(__9____1887), .CLK(clk), .Q(n520), .Q_N(n1003) );
  dfrbp_1 _______________________36183 ( .D(__9____1882), .CLK(clk), .RESET_B(
        rst), .Q(n1031), .Q_N(n531) );
  dfrbp_1 __________________36184 ( .D(__9_9__1884), .CLK(clk), .RESET_B(rst), 
        .Q(n1019) );
  dfxbp_1 ______________ ( .D(__9____1881), .CLK(clk), .Q(n999), .Q_N(n536) );
  dfxbp_1 ______________36194 ( .D(__9____1869), .CLK(clk), .Q_N(n1012) );
  dfrbp_1 _______________________36195 ( .D(__9____1860), .CLK(clk), .RESET_B(
        rst), .Q(n1029), .Q_N(n535) );
  dfxbp_1 ____________0_ ( .D(__9_9), .CLK(clk), .Q(n1011), .Q_N(n537) );
  dfxbp_1 ______________36198 ( .D(__9____1861), .CLK(clk), .Q(n1013), .Q_N(
        n533) );
  dfxbp_1 ______________36199 ( .D(__9____1872), .CLK(clk), .Q(n1007), .Q_N(
        n523) );
  dfxbp_1 ______________36200 ( .D(__9____1870), .CLK(clk), .Q_N(n1009) );
  dfxbp_1 ______________36201 ( .D(__9____1868), .CLK(clk), .Q(n534), .Q_N(
        n1010) );
  dfxbp_1 ______________36202 ( .D(__9____1873), .CLK(clk), .Q_N(n1006) );
  dfrbp_1 __________________36209 ( .D(__90___1854), .CLK(clk), .RESET_B(rst), 
        .Q(n530), .Q_N(n1025) );
  dfrbp_1 _______________________36221 ( .D(__90_), .CLK(clk), .RESET_B(rst), 
        .Q(n529), .Q_N(n1000) );
  dfrbp_1 __________________36229 ( .D(___99__1850), .CLK(clk), .RESET_B(rst), 
        .Q(n516), .Q_N(n1021) );
  dfxbp_1 __________________36230 ( .D(____0___2025), .CLK(clk), .Q_N(n1015)
         );
  dfrbp_1 __________________36246 ( .D(_______1827), .CLK(clk), .RESET_B(rst), 
        .Q(n1024) );
  dfrbp_1 ____0__________________ ( .D(_______1830), .CLK(clk), .RESET_B(rst), 
        .Q(n525), .Q_N(n1004) );
  dfxbp_1 __________________36247 ( .D(_______1826), .CLK(clk), .Q_N(
        _______________1154) );
  dfxbp_1 __________________36250 ( .D(_______1828), .CLK(clk), .Q(n1018) );
  dfrbp_1 ____0__________________36256 ( .D(_______1820), .CLK(clk), .RESET_B(
        rst), .Q(n519), .Q_N(n1001) );
  dfxbp_1 __________________36259 ( .D(n47), .CLK(clk), .Q_N(___09___2013) );
  dfrbp_1 ____0__________________36260 ( .D(____0__1814), .CLK(clk), .RESET_B(
        rst), .Q(n526), .Q_N(n1017) );
  dfrbp_1 ____0__________________36268 ( .D(_______1806), .CLK(clk), .RESET_B(
        rst), .Q(n515), .Q_N(n1005) );
  dfrbp_1 ____0__________________36271 ( .D(_______1801), .CLK(clk), .RESET_B(
        rst), .Q(n528), .Q_N(n1032) );
  dfrbp_1 ________________0_ ( .D(_______1793), .CLK(clk), .RESET_B(rst), .Q(
        n1022), .Q_N(n524) );
  dfrbp_1 _____________________0_ ( .D(_______1798), .CLK(clk), .RESET_B(rst), 
        .Q_N(n1030) );
  dfrbp_1 ____0__________________36274 ( .D(_______1794), .CLK(clk), .RESET_B(
        rst), .Q(n521), .Q_N(n1033) );
  dfxbp_1 __________________36279 ( .D(n48), .CLK(clk), .Q(n159), .Q_N(valid)
         );
  dfrbp_1 ____0________________0_ ( .D(_______1781), .CLK(clk), .RESET_B(rst), 
        .Q(n514), .Q_N(n1028) );
  dfxbp_1 ________________0_36303 ( .D(___0___1764), .CLK(clk), .Q(
        ___________0___1152) );
  dfrbp_1 ____0__________________36334 ( .D(n2), .CLK(clk), .RESET_B(rst), .Q(
        n527), .Q_N(n1002) );
  dfrbp_1 ____0________________0_36396 ( .D(_______1652), .CLK(clk), .RESET_B(
        rst), .Q(n518), .Q_N(n1008) );
  dfrbp_1 __________________36586 ( .D(_______1397), .CLK(clk), .RESET_B(rst), 
        .Q(n1026) );
  inv_1 U527 ( .A(n540), .Y(n48) );
  inv_1 U528 ( .A(n541), .Y(n47) );
  a21oi_1 U529 ( .A1(n542), .A2(n543), .B1(n1030), .Y(n541) );
  nand2_1 U530 ( .A(n544), .B(n545), .Y(n45) );
  mux2_1 U531 ( .A0(n1015), .A1(n546), .S(n547), .X(n544) );
  a21oi_1 U532 ( .A1(n1026), .A2(n1016), .B1(n548), .Y(n546) );
  nand4_1 U533 ( .A(n549), .B(n550), .C(n551), .D(n552), .Y(n2) );
  inv_1 U534 ( .A(_______1652), .Y(n552) );
  or3_1 U535 ( .A(n553), .B(n515), .C(n554), .X(n550) );
  nand3_1 U536 ( .A(n555), .B(n556), .C(n557), .Y(n549) );
  o221ai_1 U537 ( .A1(n553), .A2(n558), .B1(n1004), .B2(n559), .C1(n560), .Y(
        _______1830) );
  nor3_1 U538 ( .A(n561), .B(n562), .C(n563), .Y(n560) );
  inv_1 U539 ( .A(n564), .Y(n562) );
  nor3_1 U540 ( .A(n565), .B(n1001), .C(n566), .Y(n561) );
  o21ai_0 U541 ( .A1(n567), .A2(n568), .B1(n569), .Y(n558) );
  o22ai_1 U542 ( .A1(n515), .A2(n554), .B1(n570), .B2(n525), .Y(n569) );
  nor4_1 U543 ( .A(n571), .B(n572), .C(n573), .D(n574), .Y(n570) );
  inv_1 U544 ( .A(n575), .Y(n572) );
  nor3_1 U545 ( .A(n576), .B(n577), .C(n578), .Y(n567) );
  nand3_1 U546 ( .A(datain[7]), .B(n579), .C(datain[0]), .Y(n576) );
  mux2i_1 U547 ( .A0(n580), .A1(n581), .S(n582), .Y(_______1828) );
  a21oi_1 U548 ( .A1(n583), .A2(n520), .B1(n584), .Y(n581) );
  nand3_1 U549 ( .A(n1020), .B(n585), .C(clk), .Y(n580) );
  nor2_1 U550 ( .A(n586), .B(n159), .Y(_______1827) );
  nor2_1 U551 ( .A(n587), .B(n586), .Y(_______1826) );
  inv_1 U552 ( .A(n588), .Y(n586) );
  o211ai_1 U553 ( .A1(n566), .A2(n565), .B1(n589), .C1(n590), .Y(_______1820)
         );
  a21oi_1 U554 ( .A1(n1001), .A2(n591), .B1(n563), .Y(n590) );
  inv_1 U555 ( .A(n592), .Y(n563) );
  o211ai_1 U556 ( .A1(n1001), .A2(n593), .B1(n594), .C1(n595), .Y(n592) );
  nor4_1 U557 ( .A(op[0]), .B(n577), .C(n596), .D(n597), .Y(n593) );
  o221ai_1 U558 ( .A1(n598), .A2(n565), .B1(n527), .B2(n599), .C1(n600), .Y(
        n591) );
  or4_1 U559 ( .A(n601), .B(n573), .C(n602), .D(n603), .X(n600) );
  a21oi_1 U560 ( .A1(n1005), .A2(n554), .B1(n1004), .Y(n598) );
  nand4_1 U561 ( .A(n604), .B(n605), .C(n575), .D(n577), .Y(n554) );
  mux2i_1 U562 ( .A0(n606), .A1(n607), .S(n525), .Y(n589) );
  nor3_1 U563 ( .A(n608), .B(op[0]), .C(n559), .Y(n606) );
  inv_1 U564 ( .A(n555), .Y(n565) );
  inv_1 U565 ( .A(n609), .Y(n566) );
  o22ai_1 U566 ( .A1(n610), .A2(n568), .B1(datain[5]), .B2(n611), .Y(n609) );
  mux2i_1 U567 ( .A0(n612), .A1(n613), .S(n515), .Y(n611) );
  nor2_1 U568 ( .A(n579), .B(n614), .Y(n613) );
  mux2i_1 U569 ( .A0(n615), .A1(n616), .S(n525), .Y(n614) );
  nor3_1 U570 ( .A(n617), .B(n618), .C(n619), .Y(n616) );
  nand3_1 U571 ( .A(n620), .B(n519), .C(n621), .Y(n617) );
  nor3_1 U572 ( .A(n596), .B(n620), .C(n602), .Y(n615) );
  nor3_1 U573 ( .A(n597), .B(n622), .C(n596), .Y(n612) );
  nand4_1 U574 ( .A(n623), .B(n564), .C(n551), .D(n624), .Y(_______1806) );
  inv_1 U575 ( .A(n607), .Y(n624) );
  a21oi_1 U576 ( .A1(n622), .A2(n625), .B1(n559), .Y(n607) );
  nand4_1 U577 ( .A(n1008), .B(n515), .C(n527), .D(n519), .Y(n559) );
  or2_0 U578 ( .A(n553), .B(n568), .X(n551) );
  inv_1 U579 ( .A(n557), .Y(n568) );
  nand2_1 U580 ( .A(n1001), .B(n555), .Y(n553) );
  nand4_1 U581 ( .A(n518), .B(n527), .C(n626), .D(n627), .Y(n564) );
  a21oi_1 U582 ( .A1(n525), .A2(n519), .B1(n628), .Y(n627) );
  mux2i_1 U583 ( .A0(n519), .A1(n525), .S(n515), .Y(n628) );
  nand3_1 U584 ( .A(datain[1]), .B(n620), .C(n629), .Y(n626) );
  mux2i_1 U585 ( .A0(n630), .A1(n631), .S(n519), .Y(n629) );
  nand3_1 U586 ( .A(datain[5]), .B(n621), .C(n632), .Y(n631) );
  or3_1 U587 ( .A(n618), .B(datain[5]), .C(n633), .X(n630) );
  nand3_1 U588 ( .A(n557), .B(n555), .C(n610), .Y(n623) );
  inv_1 U589 ( .A(n556), .Y(n610) );
  nand3_1 U590 ( .A(n634), .B(n604), .C(n635), .Y(n556) );
  nor3_1 U591 ( .A(n577), .B(datain[7]), .C(n579), .Y(n635) );
  nor2_1 U592 ( .A(n527), .B(n518), .Y(n555) );
  o211ai_1 U593 ( .A1(n1032), .A2(n636), .B1(n637), .C1(n638), .Y(_______1801)
         );
  mux2i_1 U594 ( .A0(n639), .A1(n640), .S(n514), .Y(n638) );
  o221ai_1 U595 ( .A1(n641), .A2(n642), .B1(n643), .B2(n644), .C1(n645), .Y(
        n640) );
  nand2_1 U596 ( .A(n646), .B(n647), .Y(n642) );
  inv_1 U597 ( .A(n648), .Y(n639) );
  a221oi_1 U598 ( .A1(n649), .A2(n650), .B1(n651), .B2(n646), .C1(n652), .Y(
        n648) );
  o211ai_1 U599 ( .A1(n653), .A2(n644), .B1(n654), .C1(n655), .Y(n652) );
  or3_1 U600 ( .A(n656), .B(n657), .C(n658), .X(n655) );
  inv_1 U601 ( .A(n659), .Y(n637) );
  nand4_1 U602 ( .A(n660), .B(n661), .C(n662), .D(n663), .Y(_______1798) );
  nor4_1 U603 ( .A(n664), .B(n665), .C(n666), .D(n667), .Y(n663) );
  inv_1 U604 ( .A(n668), .Y(n664) );
  nor2_1 U605 ( .A(n669), .B(n670), .Y(n662) );
  nand4_1 U606 ( .A(n671), .B(n672), .C(n673), .D(n520), .Y(n661) );
  o221ai_1 U607 ( .A1(n674), .A2(n675), .B1(n1032), .B2(n676), .C1(n677), .Y(
        _______1794) );
  o21ai_0 U608 ( .A1(n678), .A2(n679), .B1(n646), .Y(n677) );
  mux2i_1 U609 ( .A0(n680), .A1(n514), .S(n528), .Y(n679) );
  nand2_1 U610 ( .A(n681), .B(n514), .Y(n680) );
  nor2_1 U611 ( .A(n682), .B(n683), .Y(n676) );
  inv_1 U612 ( .A(n636), .Y(n683) );
  nand3_1 U613 ( .A(n521), .B(n514), .C(n684), .Y(n636) );
  o32ai_1 U614 ( .A1(n685), .A2(n608), .A3(n658), .B1(n686), .B2(n687), .Y(
        n684) );
  mux2i_1 U615 ( .A0(n651), .A1(n688), .S(n514), .Y(n675) );
  nor2_1 U616 ( .A(n689), .B(n690), .Y(n688) );
  inv_1 U617 ( .A(n678), .Y(n690) );
  nand2_1 U618 ( .A(n588), .B(___________0___1152), .Y(_______1793) );
  nand4_1 U619 ( .A(n691), .B(n692), .C(n693), .D(n694), .Y(_______1781) );
  a221oi_1 U620 ( .A1(n682), .A2(n647), .B1(n695), .B2(n678), .C1(n659), .Y(
        n694) );
  nand2_1 U621 ( .A(n696), .B(n697), .Y(n659) );
  nand4_1 U622 ( .A(n698), .B(n678), .C(n699), .D(n700), .Y(n697) );
  nor3_1 U623 ( .A(n597), .B(n514), .C(n577), .Y(n700) );
  nand4_1 U624 ( .A(n701), .B(n649), .C(n647), .D(n702), .Y(n696) );
  and3_1 U625 ( .A(n1028), .B(n656), .C(n698), .X(n682) );
  nand4_1 U626 ( .A(n703), .B(datain[2]), .C(datain[5]), .D(n704), .Y(n656) );
  nand2_1 U627 ( .A(n705), .B(n706), .Y(n693) );
  mux2i_1 U628 ( .A0(n707), .A1(n708), .S(n514), .Y(n705) );
  nor2_1 U629 ( .A(n608), .B(n685), .Y(n708) );
  nand3_1 U630 ( .A(n709), .B(n514), .C(n646), .Y(n691) );
  o21ai_0 U631 ( .A1(n1032), .A2(n710), .B1(n657), .Y(n709) );
  inv_1 U632 ( .A(n647), .Y(n657) );
  o221ai_1 U633 ( .A1(n519), .A2(n599), .B1(n702), .B2(n594), .C1(n601), .Y(
        _______1652) );
  nand3_1 U634 ( .A(n518), .B(n527), .C(n557), .Y(n601) );
  nor2_1 U635 ( .A(n525), .B(n515), .Y(n557) );
  nand4_1 U636 ( .A(datain[5]), .B(datain[0]), .C(n704), .D(n621), .Y(n594) );
  nand3_1 U637 ( .A(n515), .B(n525), .C(n518), .Y(n599) );
  nand2_1 U638 ( .A(n545), .B(n538), .Y(_______1397) );
  nand2_1 U639 ( .A(n711), .B(n545), .Y(____0___2025) );
  mux2i_1 U640 ( .A0(n712), .A1(n713), .S(n547), .Y(n711) );
  nand2_1 U641 ( .A(op[0]), .B(n714), .Y(n713) );
  xor2_1 U642 ( .A(n1023), .B(n548), .X(n714) );
  a21oi_1 U643 ( .A1(n715), .A2(n1014), .B1(n584), .Y(n712) );
  nor2_1 U644 ( .A(n1003), .B(n716), .Y(n715) );
  nand3_1 U645 ( .A(n717), .B(n654), .C(n718), .Y(____0__1814) );
  a21oi_1 U646 ( .A1(n695), .A2(n1032), .B1(n719), .Y(n718) );
  mux2i_1 U647 ( .A0(n720), .A1(n721), .S(n514), .Y(n719) );
  nor4_1 U648 ( .A(n722), .B(n723), .C(n724), .D(n706), .Y(n721) );
  inv_1 U649 ( .A(n645), .Y(n724) );
  nand3_1 U650 ( .A(n698), .B(n678), .C(n689), .Y(n645) );
  and3_1 U651 ( .A(n725), .B(n575), .C(n726), .X(n689) );
  nor3_1 U652 ( .A(n727), .B(n728), .C(n577), .Y(n726) );
  nor2_1 U653 ( .A(n528), .B(n1033), .Y(n678) );
  nor3_1 U654 ( .A(n687), .B(n710), .C(n729), .Y(n723) );
  inv_1 U655 ( .A(n686), .Y(n710) );
  nand2_1 U656 ( .A(n730), .B(datain[5]), .Y(n686) );
  o22ai_1 U657 ( .A1(n731), .A2(n692), .B1(n681), .B2(n644), .Y(n722) );
  inv_1 U658 ( .A(n732), .Y(n644) );
  inv_1 U659 ( .A(n643), .Y(n681) );
  nand2_1 U660 ( .A(n730), .B(n577), .Y(n643) );
  and3_1 U661 ( .A(n733), .B(n734), .C(n735), .X(n730) );
  nor3_1 U662 ( .A(n727), .B(datain[1]), .C(n620), .Y(n735) );
  inv_1 U663 ( .A(n650), .Y(n692) );
  nor4_1 U664 ( .A(n736), .B(n737), .C(n573), .D(n738), .Y(n731) );
  nand3_1 U665 ( .A(datain[1]), .B(n620), .C(datain[2]), .Y(n736) );
  a222oi_1 U666 ( .A1(n647), .A2(n702), .B1(n732), .B2(n653), .C1(n650), .C2(
        n739), .Y(n720) );
  inv_1 U667 ( .A(n649), .Y(n739) );
  nor3_1 U668 ( .A(datain[6]), .B(op[1]), .C(n608), .Y(n649) );
  inv_1 U669 ( .A(n625), .Y(n608) );
  nor3_1 U670 ( .A(n573), .B(n597), .C(n738), .Y(n625) );
  nand2_1 U671 ( .A(n618), .B(n577), .Y(n573) );
  nor2_1 U672 ( .A(n658), .B(n740), .Y(n650) );
  nand4_1 U673 ( .A(n741), .B(datain[7]), .C(n703), .D(n742), .Y(n653) );
  nor3_1 U674 ( .A(n579), .B(datain[5]), .C(datain[2]), .Y(n742) );
  nor2_1 U675 ( .A(n687), .B(n740), .Y(n732) );
  inv_1 U676 ( .A(n646), .Y(n687) );
  and4_1 U677 ( .A(n701), .B(n734), .C(n725), .D(n743), .X(n695) );
  nor3_1 U678 ( .A(n597), .B(n674), .C(n577), .Y(n743) );
  nand2_1 U679 ( .A(n575), .B(n727), .Y(n597) );
  nor2_1 U680 ( .A(datain[7]), .B(datain[1]), .Y(n575) );
  nand2_1 U681 ( .A(n706), .B(n707), .Y(n654) );
  nor2_1 U682 ( .A(n658), .B(n729), .Y(n706) );
  inv_1 U683 ( .A(n698), .Y(n658) );
  nor2_1 U684 ( .A(n1017), .B(n674), .Y(n698) );
  nand3_1 U685 ( .A(n647), .B(n641), .C(n646), .Y(n717) );
  nor2_1 U686 ( .A(n526), .B(n674), .Y(n646) );
  inv_1 U687 ( .A(n702), .Y(n674) );
  nand2_1 U688 ( .A(n595), .B(n1001), .Y(n702) );
  nor4_1 U689 ( .A(n515), .B(n518), .C(n1004), .D(n1002), .Y(n595) );
  nand4_1 U690 ( .A(n727), .B(n577), .C(n704), .D(n744), .Y(n641) );
  nor2_1 U691 ( .A(n618), .B(n685), .Y(n744) );
  inv_1 U692 ( .A(n603), .Y(n704) );
  nand3_1 U693 ( .A(datain[1]), .B(n745), .C(datain[7]), .Y(n603) );
  mux2i_1 U694 ( .A0(___09___2013), .A1(n746), .S(n747), .Y(___99__1850) );
  nor3_1 U695 ( .A(n748), .B(n749), .C(n750), .Y(n746) );
  mux2i_1 U696 ( .A0(n751), .A1(n530), .S(n516), .Y(n748) );
  nand2_1 U697 ( .A(n530), .B(n520), .Y(n751) );
  nor2_1 U698 ( .A(n542), .B(___0____2003), .Y(___0____1999) );
  nor2_1 U699 ( .A(n542), .B(___0____2004), .Y(___0____1998) );
  nor2_1 U700 ( .A(n542), .B(___0____2008), .Y(___0____1997) );
  nand2_1 U701 ( .A(n540), .B(n124), .Y(___0____1994) );
  nor2_1 U702 ( .A(n542), .B(___0____2005), .Y(___0____1992) );
  nor2_1 U703 ( .A(n542), .B(___0____2006), .Y(___0____1991) );
  o211ai_1 U704 ( .A1(n1012), .A2(n752), .B1(n753), .C1(n754), .Y(___0____1990) );
  xnor2_1 U705 ( .A(n755), .B(n518), .Y(n754) );
  nand3_1 U706 ( .A(n1019), .B(n756), .C(n757), .Y(n755) );
  o221ai_1 U707 ( .A1(n758), .A2(n759), .B1(n537), .B2(n752), .C1(n760), .Y(
        ___0____1989) );
  inv_1 U708 ( .A(n761), .Y(n758) );
  o21ai_0 U709 ( .A1(n1012), .A2(n1011), .B1(n762), .Y(n761) );
  o221ai_1 U710 ( .A1(n759), .A2(n763), .B1(n533), .B2(n752), .C1(n760), .Y(
        ___0____1987) );
  or2_0 U711 ( .A(n764), .B(n765), .X(n760) );
  xnor2_1 U712 ( .A(n766), .B(n767), .Y(n763) );
  xnor2_1 U713 ( .A(n1009), .B(n768), .Y(n767) );
  o21ai_0 U714 ( .A1(n1006), .A2(n752), .B1(n769), .Y(___0____1985) );
  o21ai_0 U715 ( .A1(n523), .A2(n752), .B1(n769), .Y(___0____1983) );
  inv_1 U716 ( .A(n770), .Y(n769) );
  o221ai_1 U717 ( .A1(n759), .A2(n771), .B1(n1010), .B2(n752), .C1(n764), .Y(
        ___0____1982) );
  xor2_1 U718 ( .A(n772), .B(n773), .X(n771) );
  xnor2_1 U719 ( .A(n774), .B(n775), .Y(n773) );
  xnor2_1 U720 ( .A(n1006), .B(n518), .Y(n772) );
  o221ai_1 U721 ( .A1(n759), .A2(n776), .B1(n536), .B2(n752), .C1(n764), .Y(
        ___0____1981) );
  nand2_1 U722 ( .A(n777), .B(n778), .Y(n764) );
  xor2_1 U723 ( .A(n779), .B(n780), .X(n776) );
  xnor2_1 U724 ( .A(n781), .B(n1007), .Y(n780) );
  nand2_1 U725 ( .A(n588), .B(n782), .Y(___0___1764) );
  nand3_1 U726 ( .A(n783), .B(n516), .C(n1022), .Y(n782) );
  a21oi_1 U727 ( .A1(n784), .A2(n647), .B1(n785), .Y(n588) );
  mux2_1 U728 ( .A0(n786), .A1(n651), .S(n1028), .X(n785) );
  nor2_1 U729 ( .A(n740), .B(n526), .Y(n786) );
  nor2_1 U730 ( .A(n521), .B(n1032), .Y(n647) );
  nand2_1 U731 ( .A(n540), .B(n125), .Y(___0_9__1995) );
  nor2_1 U732 ( .A(n542), .B(n1030), .Y(n540) );
  nor2_1 U733 ( .A(n542), .B(___0____2007), .Y(___0_0__1996) );
  o21ai_0 U734 ( .A1(n1009), .A2(n752), .B1(n753), .Y(___09___2017) );
  a21oi_1 U735 ( .A1(n777), .A2(n765), .B1(n770), .Y(n753) );
  o22ai_1 U736 ( .A1(n778), .A2(n787), .B1(n788), .B2(n756), .Y(n770) );
  o22ai_1 U737 ( .A1(n781), .A2(n779), .B1(n789), .B2(n523), .Y(n756) );
  and2_0 U738 ( .A(n779), .B(n781), .X(n789) );
  xnor2_1 U739 ( .A(n999), .B(n790), .Y(n779) );
  inv_1 U740 ( .A(n791), .Y(n781) );
  o22ai_1 U741 ( .A1(n774), .A2(n792), .B1(n1006), .B2(n793), .Y(n791) );
  nor2_1 U742 ( .A(n775), .B(n794), .Y(n793) );
  inv_1 U743 ( .A(n775), .Y(n792) );
  xnor2_1 U744 ( .A(n1010), .B(n790), .Y(n775) );
  inv_1 U745 ( .A(n794), .Y(n774) );
  o22ai_1 U746 ( .A1(n766), .A2(n768), .B1(n1009), .B2(n795), .Y(n794) );
  and2_0 U747 ( .A(n768), .B(n766), .X(n795) );
  o21ai_0 U748 ( .A1(n1011), .A2(n790), .B1(n762), .Y(n768) );
  xnor2_1 U749 ( .A(n533), .B(n788), .Y(n766) );
  inv_1 U750 ( .A(n790), .Y(n788) );
  nor2_1 U751 ( .A(n759), .B(n1019), .Y(n790) );
  xnor2_1 U752 ( .A(n796), .B(n1008), .Y(n778) );
  o22ai_1 U753 ( .A1(n523), .A2(n797), .B1(n999), .B2(n798), .Y(n796) );
  nor2_1 U754 ( .A(n799), .B(n1007), .Y(n798) );
  inv_1 U755 ( .A(n799), .Y(n797) );
  a21oi_1 U756 ( .A1(n534), .A2(n800), .B1(n801), .Y(n799) );
  xnor2_1 U757 ( .A(n802), .B(n1008), .Y(n801) );
  o21ai_0 U758 ( .A1(n534), .A2(n800), .B1(n1006), .Y(n802) );
  nand2_1 U759 ( .A(n803), .B(n804), .Y(n800) );
  o22ai_1 U760 ( .A1(n1011), .A2(n1012), .B1(n1009), .B2(n1013), .Y(n803) );
  and3_1 U761 ( .A(n762), .B(n804), .C(n805), .X(n765) );
  a22oi_1 U762 ( .A1(n1006), .A2(n534), .B1(n999), .B2(n523), .Y(n805) );
  nand2_1 U763 ( .A(n1009), .B(n1013), .Y(n804) );
  nand2_1 U764 ( .A(n1011), .B(n1012), .Y(n762) );
  mux2i_1 U765 ( .A0(n806), .A1(n807), .S(n747), .Y(__9____1926) );
  a211oi_1 U766 ( .A1(n530), .A2(n520), .B1(n750), .C1(n622), .Y(n807) );
  o211ai_1 U767 ( .A1(n530), .A2(n520), .B1(n1017), .C1(n651), .Y(n750) );
  nor3_1 U768 ( .A(n524), .B(n583), .C(n808), .Y(n806) );
  mux2i_1 U769 ( .A0(n809), .A1(n539), .S(n582), .Y(__9____1920) );
  nor2_1 U770 ( .A(n810), .B(n811), .Y(n809) );
  xor2_1 U771 ( .A(n812), .B(n1014), .X(n811) );
  nand2_1 U772 ( .A(n813), .B(n814), .Y(__9____1911) );
  nor4_1 U773 ( .A(n815), .B(n816), .C(n817), .D(n818), .Y(n814) );
  a21oi_1 U774 ( .A1(n819), .A2(n634), .B1(n820), .Y(n818) );
  a21oi_1 U775 ( .A1(n821), .A2(n734), .B1(n822), .Y(n817) );
  a21oi_1 U776 ( .A1(n823), .A2(n824), .B1(n825), .Y(n816) );
  nand4_1 U777 ( .A(n826), .B(n668), .C(n827), .D(n828), .Y(n815) );
  nand3_1 U778 ( .A(n829), .B(n604), .C(n670), .Y(n826) );
  nor4_1 U779 ( .A(n830), .B(n831), .C(n832), .D(n833), .Y(n813) );
  o221ai_1 U780 ( .A1(n834), .A2(n835), .B1(n836), .B2(n837), .C1(n838), .Y(
        n830) );
  inv_1 U781 ( .A(n839), .Y(n836) );
  a222oi_1 U782 ( .A1(n840), .A2(n841), .B1(n842), .B2(n671), .C1(n843), .C2(
        n844), .Y(n834) );
  nand3_1 U783 ( .A(n634), .B(n741), .C(n845), .Y(n844) );
  inv_1 U784 ( .A(n846), .Y(n840) );
  nand4_1 U785 ( .A(n847), .B(n848), .C(n849), .D(n850), .Y(__9____1899) );
  nor4_1 U786 ( .A(n851), .B(n852), .C(n853), .D(n854), .Y(n850) );
  o22ai_1 U787 ( .A1(n855), .A2(n856), .B1(n857), .B2(n858), .Y(n852) );
  inv_1 U788 ( .A(n859), .Y(n857) );
  a221oi_1 U789 ( .A1(n860), .A2(n671), .B1(n861), .B2(n862), .C1(n863), .Y(
        n855) );
  o21ai_0 U790 ( .A1(n864), .A2(n865), .B1(n824), .Y(n863) );
  inv_1 U791 ( .A(n838), .Y(n851) );
  nor4_1 U792 ( .A(n866), .B(n667), .C(n669), .D(n867), .Y(n838) );
  o32ai_1 U793 ( .A1(n837), .A2(n868), .A3(n869), .B1(n870), .B2(n871), .Y(
        n867) );
  nand2_1 U794 ( .A(n666), .B(n632), .Y(n871) );
  inv_1 U795 ( .A(n872), .Y(n866) );
  and3_1 U796 ( .A(n873), .B(n822), .C(n874), .X(n849) );
  o21ai_0 U797 ( .A1(n875), .A2(n876), .B1(n841), .Y(n848) );
  and3_1 U798 ( .A(n877), .B(n745), .C(n672), .X(n875) );
  o21ai_0 U799 ( .A1(n878), .A2(n879), .B1(n861), .Y(n847) );
  a21oi_1 U800 ( .A1(n877), .A2(n880), .B1(n825), .Y(n878) );
  o32ai_1 U801 ( .A1(n881), .A2(n747), .A3(n808), .B1(n882), .B2(n883), .Y(
        __9____1887) );
  nand2_1 U802 ( .A(n1021), .B(op[0]), .Y(n883) );
  nand4_1 U803 ( .A(n884), .B(n660), .C(n885), .D(n886), .Y(__9____1882) );
  and4_1 U804 ( .A(n887), .B(n872), .C(n888), .D(n889), .X(n886) );
  a222oi_1 U805 ( .A1(n890), .A2(n891), .B1(n876), .B2(n892), .C1(n893), .C2(
        n894), .Y(n889) );
  o21ai_0 U806 ( .A1(n842), .A2(n895), .B1(n896), .Y(n892) );
  nor3_1 U807 ( .A(n574), .B(n897), .C(n685), .Y(n842) );
  o221ai_1 U808 ( .A1(n898), .A2(n864), .B1(n824), .B2(n899), .C1(n823), .Y(
        n891) );
  o21ai_0 U809 ( .A1(n897), .A2(n870), .B1(n670), .Y(n888) );
  inv_1 U810 ( .A(n900), .Y(n670) );
  inv_1 U811 ( .A(n604), .Y(n897) );
  nor2_1 U812 ( .A(n571), .B(n618), .Y(n604) );
  nand3_1 U813 ( .A(n901), .B(n880), .C(n667), .Y(n887) );
  inv_1 U814 ( .A(n902), .Y(n667) );
  a222oi_1 U815 ( .A1(n669), .A2(n846), .B1(n672), .B2(n903), .C1(n879), .C2(
        n839), .Y(n885) );
  nand2_1 U816 ( .A(n896), .B(n904), .Y(n839) );
  nand3_1 U817 ( .A(n699), .B(n621), .C(n905), .Y(n904) );
  inv_1 U818 ( .A(n906), .Y(n669) );
  and3_1 U819 ( .A(n907), .B(n908), .C(n822), .X(n660) );
  inv_1 U820 ( .A(n909), .Y(n884) );
  nor2_1 U821 ( .A(n808), .B(n910), .Y(__9____1881) );
  nor2_1 U822 ( .A(n808), .B(n911), .Y(__9____1873) );
  nor2_1 U823 ( .A(n808), .B(n620), .Y(__9____1872) );
  inv_1 U824 ( .A(datain[7]), .Y(n620) );
  nor2_1 U825 ( .A(n808), .B(n577), .Y(__9____1870) );
  inv_1 U826 ( .A(datain[5]), .Y(n577) );
  nor2_1 U827 ( .A(n808), .B(n749), .Y(__9____1869) );
  nor2_1 U828 ( .A(n808), .B(n727), .Y(__9____1868) );
  nor2_1 U829 ( .A(n808), .B(n579), .Y(__9____1861) );
  inv_1 U830 ( .A(datain[1]), .Y(n579) );
  nand3_1 U831 ( .A(n912), .B(n913), .C(n914), .Y(__9____1860) );
  nor4_1 U832 ( .A(n915), .B(n916), .C(n666), .D(n917), .Y(n914) );
  nor3_1 U833 ( .A(n918), .B(n869), .C(n835), .Y(n917) );
  inv_1 U834 ( .A(n919), .Y(n869) );
  o32ai_1 U835 ( .A1(n837), .A2(n898), .A3(n823), .B1(n920), .B2(n921), .Y(
        n916) );
  nand2_1 U836 ( .A(n741), .B(n922), .Y(n921) );
  o32ai_1 U837 ( .A1(n835), .A2(n896), .A3(n923), .B1(n924), .B2(n820), .Y(
        n922) );
  inv_1 U838 ( .A(n843), .Y(n896) );
  inv_1 U839 ( .A(n861), .Y(n823) );
  inv_1 U840 ( .A(n865), .Y(n898) );
  nand2_1 U841 ( .A(n821), .B(n741), .Y(n865) );
  nand4_1 U842 ( .A(n925), .B(n907), .C(n872), .D(n828), .Y(n915) );
  nand3_1 U843 ( .A(n890), .B(n861), .C(n926), .Y(n828) );
  nand3_1 U844 ( .A(n672), .B(n919), .C(n868), .Y(n872) );
  nand2_1 U845 ( .A(n927), .B(n928), .Y(n907) );
  nor3_1 U846 ( .A(n929), .B(n930), .C(n931), .Y(n913) );
  a21oi_1 U847 ( .A1(n901), .A2(n880), .B1(n902), .Y(n931) );
  nand4_1 U848 ( .A(n1029), .B(n843), .C(n932), .D(n531), .Y(n902) );
  inv_1 U849 ( .A(n933), .Y(n930) );
  o21ai_0 U850 ( .A1(n923), .A2(n602), .B1(n854), .Y(n933) );
  nand2_1 U851 ( .A(n934), .B(n908), .Y(n854) );
  o22ai_1 U852 ( .A1(n745), .A2(n934), .B1(n846), .B2(n906), .Y(n929) );
  nand2_1 U853 ( .A(n905), .B(n935), .Y(n906) );
  nor4_1 U854 ( .A(n832), .B(n853), .C(n936), .D(n937), .Y(n912) );
  mux2i_1 U855 ( .A0(n938), .A1(n908), .S(n738), .Y(n937) );
  inv_1 U856 ( .A(n734), .Y(n738) );
  nand2_1 U857 ( .A(n939), .B(n821), .Y(n938) );
  inv_1 U858 ( .A(n822), .Y(n939) );
  nand4_1 U859 ( .A(n905), .B(n1029), .C(n932), .D(n531), .Y(n822) );
  o21ai_0 U860 ( .A1(n940), .A2(n894), .B1(n900), .Y(n853) );
  nand4_1 U861 ( .A(n919), .B(n1029), .C(n1031), .D(n932), .Y(n900) );
  nand2_1 U862 ( .A(n941), .B(n734), .Y(n894) );
  o32ai_1 U863 ( .A1(n856), .A2(n860), .A3(n895), .B1(n859), .B2(n858), .Y(
        n832) );
  nand3_1 U864 ( .A(n734), .B(n942), .C(n725), .Y(n859) );
  o22ai_1 U865 ( .A1(n582), .A2(n943), .B1(n1018), .B2(n944), .Y(__9_9__1884)
         );
  nor2_1 U866 ( .A(n582), .B(n532), .Y(n944) );
  and3_1 U867 ( .A(op[0]), .B(n812), .C(n585), .X(n943) );
  nor2_1 U868 ( .A(n808), .B(n618), .Y(__9_9) );
  inv_1 U869 ( .A(n945), .Y(n808) );
  nand2_1 U870 ( .A(n946), .B(n545), .Y(__99___1933) );
  mux2i_1 U871 ( .A0(n947), .A1(n948), .S(n547), .Y(n946) );
  nor2_1 U872 ( .A(n949), .B(n701), .Y(n547) );
  a21oi_1 U873 ( .A1(n514), .A2(n950), .B1(n951), .Y(n949) );
  o21ai_0 U874 ( .A1(n526), .A2(n1032), .B1(n521), .Y(n950) );
  xnor2_1 U875 ( .A(n1015), .B(n548), .Y(n948) );
  nor2_1 U876 ( .A(n1016), .B(n1026), .Y(n548) );
  a21oi_1 U877 ( .A1(n583), .A2(n952), .B1(n584), .Y(n947) );
  or2_0 U878 ( .A(n520), .B(n1014), .X(n952) );
  nor2_1 U879 ( .A(n622), .B(n953), .Y(__99___1932) );
  mux2i_1 U880 ( .A0(n954), .A1(n945), .S(n582), .Y(n953) );
  and2_0 U881 ( .A(n545), .B(n729), .X(n582) );
  mux2i_1 U882 ( .A0(n955), .A1(n951), .S(n514), .Y(n545) );
  nor2_1 U883 ( .A(n1017), .B(n1033), .Y(n955) );
  nand4_1 U884 ( .A(n752), .B(n543), .C(n759), .D(n956), .Y(n945) );
  and2_0 U885 ( .A(n787), .B(n587), .X(n956) );
  nor2_1 U886 ( .A(n584), .B(n583), .Y(n587) );
  inv_1 U887 ( .A(n716), .Y(n583) );
  nand4_1 U888 ( .A(n1021), .B(n1022), .C(n783), .D(n532), .Y(n716) );
  inv_1 U889 ( .A(n542), .Y(n584) );
  nand4_1 U890 ( .A(n1020), .B(n1022), .C(n783), .D(n516), .Y(n542) );
  inv_1 U891 ( .A(n777), .Y(n787) );
  nor4_1 U892 ( .A(n1024), .B(n1019), .C(n1026), .D(n957), .Y(n777) );
  nand2_1 U893 ( .A(n1023), .B(n958), .Y(n957) );
  inv_1 U894 ( .A(n757), .Y(n759) );
  nor2_1 U895 ( .A(n959), .B(n1026), .Y(n757) );
  inv_1 U896 ( .A(n960), .Y(n959) );
  nand4_1 U897 ( .A(n783), .B(n524), .C(n516), .D(n532), .Y(n543) );
  and4_1 U898 ( .A(n1019), .B(n1025), .C(n961), .D(n1026), .X(n783) );
  nor2_1 U899 ( .A(n1023), .B(n1024), .Y(n961) );
  nand3_1 U900 ( .A(n1019), .B(n1026), .C(n960), .Y(n752) );
  nor3_1 U901 ( .A(n1024), .B(n1023), .C(n962), .Y(n960) );
  inv_1 U902 ( .A(n958), .Y(n962) );
  nor4_1 U903 ( .A(n524), .B(n1025), .C(n1021), .D(n1020), .Y(n958) );
  nor2_1 U904 ( .A(n810), .B(n963), .Y(n954) );
  xnor2_1 U905 ( .A(n1019), .B(n812), .Y(n963) );
  nand2_1 U906 ( .A(n1018), .B(n1020), .Y(n812) );
  inv_1 U907 ( .A(n585), .Y(n810) );
  o22ai_1 U908 ( .A1(n521), .A2(n526), .B1(n1032), .B2(n964), .Y(n585) );
  nor2_1 U909 ( .A(n784), .B(n701), .Y(n964) );
  nor2_1 U910 ( .A(n526), .B(n514), .Y(n701) );
  o32ai_1 U911 ( .A1(n882), .A2(n965), .A3(n727), .B1(n747), .B2(
        _______________1154), .Y(__90___1854) );
  xnor2_1 U912 ( .A(n1027), .B(n1003), .Y(n965) );
  nand3_1 U913 ( .A(n651), .B(n1017), .C(n747), .Y(n882) );
  and2_0 U914 ( .A(n966), .B(n967), .X(n747) );
  o211ai_1 U915 ( .A1(n1028), .A2(n740), .B1(n729), .C1(n526), .Y(n967) );
  inv_1 U916 ( .A(n651), .Y(n729) );
  inv_1 U917 ( .A(n951), .Y(n740) );
  nor2_1 U918 ( .A(n528), .B(n521), .Y(n951) );
  o21ai_0 U919 ( .A1(n1032), .A2(n514), .B1(n1017), .Y(n966) );
  nand4_1 U920 ( .A(n968), .B(n969), .C(n970), .D(n971), .Y(__90_) );
  nor4_1 U921 ( .A(n972), .B(n973), .C(n665), .D(n974), .Y(n971) );
  inv_1 U922 ( .A(n858), .Y(n974) );
  nand2_1 U923 ( .A(n672), .B(n975), .Y(n858) );
  inv_1 U924 ( .A(n820), .Y(n665) );
  nand2_1 U925 ( .A(n935), .B(n975), .Y(n820) );
  nor3_1 U926 ( .A(n934), .B(n633), .C(n923), .Y(n973) );
  nand2_1 U927 ( .A(n890), .B(n905), .Y(n934) );
  nor3_1 U928 ( .A(n522), .B(n517), .C(n529), .Y(n905) );
  nand3_1 U929 ( .A(n976), .B(n977), .C(n978), .Y(n972) );
  o21ai_0 U930 ( .A1(n596), .A2(n870), .B1(n666), .Y(n978) );
  and3_1 U931 ( .A(n932), .B(n979), .C(n841), .X(n666) );
  or3_1 U932 ( .A(n895), .B(n825), .C(n673), .X(n977) );
  nand2_1 U933 ( .A(n821), .B(n880), .Y(n673) );
  and2_0 U934 ( .A(n725), .B(n621), .X(n821) );
  and2_0 U935 ( .A(n980), .B(n911), .X(n725) );
  inv_1 U936 ( .A(datain[6]), .Y(n911) );
  nand3_1 U937 ( .A(n861), .B(n862), .C(n890), .Y(n976) );
  inv_1 U938 ( .A(n926), .Y(n862) );
  nor3_1 U939 ( .A(n633), .B(datain[0]), .C(n737), .Y(n926) );
  nand2_1 U940 ( .A(n605), .B(n745), .Y(n633) );
  nor3_1 U941 ( .A(n936), .B(n831), .C(n909), .Y(n970) );
  nand4_1 U942 ( .A(n981), .B(n982), .C(n983), .D(n873), .Y(n909) );
  nand3_1 U943 ( .A(n919), .B(n918), .C(n876), .Y(n873) );
  nand3_1 U944 ( .A(n621), .B(n745), .C(n733), .Y(n918) );
  inv_1 U945 ( .A(n984), .Y(n621) );
  nand3_1 U946 ( .A(n879), .B(n919), .C(n868), .Y(n983) );
  and2_0 U947 ( .A(n901), .B(n734), .X(n868) );
  nor3_1 U948 ( .A(n522), .B(n998), .C(n529), .Y(n919) );
  inv_1 U949 ( .A(n837), .Y(n879) );
  nand3_1 U950 ( .A(n890), .B(n671), .C(n860), .Y(n982) );
  and2_0 U951 ( .A(n699), .B(n634), .X(n860) );
  and2_0 U952 ( .A(n703), .B(n880), .X(n699) );
  nor3_1 U953 ( .A(n618), .B(datain[6]), .C(n881), .Y(n703) );
  nand3_1 U954 ( .A(n841), .B(n846), .C(n876), .Y(n981) );
  nand2_1 U955 ( .A(n819), .B(n942), .Y(n846) );
  nor2_1 U956 ( .A(n924), .B(n571), .Y(n819) );
  inv_1 U957 ( .A(n741), .Y(n571) );
  o211ai_1 U958 ( .A1(n928), .A2(n874), .B1(n940), .C1(n925), .Y(n831) );
  nand3_1 U959 ( .A(n841), .B(n899), .C(n890), .Y(n925) );
  or3_1 U960 ( .A(n574), .B(n596), .C(n737), .X(n899) );
  nand2_1 U961 ( .A(datain[6]), .B(n881), .Y(n737) );
  inv_1 U962 ( .A(n632), .Y(n596) );
  nor2_1 U963 ( .A(n619), .B(datain[0]), .Y(n632) );
  inv_1 U964 ( .A(n893), .Y(n940) );
  nor2_1 U965 ( .A(n837), .B(n895), .Y(n893) );
  inv_1 U966 ( .A(n927), .Y(n874) );
  nor2_1 U967 ( .A(n707), .B(n985), .Y(n927) );
  nand3_1 U968 ( .A(n975), .B(n979), .C(n1030), .Y(n707) );
  nor3_1 U969 ( .A(n517), .B(n1000), .C(n522), .Y(n975) );
  nor3_1 U970 ( .A(n619), .B(n602), .C(n924), .Y(n928) );
  inv_1 U971 ( .A(n605), .Y(n602) );
  inv_1 U972 ( .A(n880), .Y(n619) );
  o211ai_1 U973 ( .A1(n895), .A2(n835), .B1(n986), .C1(n827), .Y(n936) );
  nand3_1 U974 ( .A(n876), .B(n845), .C(n987), .Y(n827) );
  nor3_1 U975 ( .A(n864), .B(n728), .C(n574), .Y(n987) );
  inv_1 U976 ( .A(n942), .Y(n574) );
  nor2_1 U977 ( .A(n622), .B(n727), .Y(n942) );
  inv_1 U978 ( .A(n745), .Y(n728) );
  inv_1 U979 ( .A(n923), .Y(n845) );
  inv_1 U980 ( .A(n835), .Y(n876) );
  o21ai_0 U981 ( .A1(n988), .A2(n903), .B1(n672), .Y(n986) );
  inv_1 U982 ( .A(n825), .Y(n672) );
  nand3_1 U983 ( .A(n1029), .B(n531), .C(n989), .Y(n825) );
  nand2_1 U984 ( .A(n864), .B(n990), .Y(n903) );
  nand3_1 U985 ( .A(n861), .B(n880), .C(n877), .Y(n990) );
  nor2_1 U986 ( .A(n910), .B(datain[4]), .Y(n880) );
  a21oi_1 U987 ( .A1(n877), .A2(n745), .B1(n824), .Y(n988) );
  inv_1 U988 ( .A(n841), .Y(n824) );
  nor3_1 U989 ( .A(n517), .B(n997), .C(n529), .Y(n841) );
  nor2_1 U990 ( .A(n870), .B(n618), .Y(n877) );
  inv_1 U991 ( .A(n829), .Y(n870) );
  nor2_1 U992 ( .A(n685), .B(n984), .Y(n829) );
  nand3_1 U993 ( .A(n1031), .B(n535), .C(n989), .Y(n835) );
  inv_1 U994 ( .A(n671), .Y(n895) );
  nor3_1 U995 ( .A(n1000), .B(n998), .C(n522), .Y(n671) );
  inv_1 U996 ( .A(n833), .Y(n969) );
  o32ai_1 U997 ( .A1(n908), .A2(n578), .A3(n923), .B1(n864), .B2(n856), .Y(
        n833) );
  inv_1 U998 ( .A(n991), .Y(n864) );
  nand2_1 U999 ( .A(n980), .B(datain[6]), .Y(n923) );
  nor2_1 U1000 ( .A(n618), .B(op[1]), .Y(n980) );
  inv_1 U1001 ( .A(datain[0]), .Y(n618) );
  nand3_1 U1002 ( .A(n932), .B(n979), .C(n991), .Y(n908) );
  nor3_1 U1003 ( .A(n1000), .B(n997), .C(n517), .Y(n991) );
  a21oi_1 U1004 ( .A1(n843), .A2(n992), .B1(n993), .Y(n968) );
  a21oi_1 U1005 ( .A1(n901), .A2(n741), .B1(n668), .Y(n993) );
  nand2_1 U1006 ( .A(n861), .B(n935), .Y(n668) );
  and3_1 U1007 ( .A(n932), .B(n535), .C(n1031), .X(n935) );
  nor2_1 U1008 ( .A(n985), .B(n1030), .Y(n932) );
  inv_1 U1009 ( .A(n994), .Y(n985) );
  nor3_1 U1010 ( .A(n998), .B(n997), .C(n529), .Y(n861) );
  nor2_1 U1011 ( .A(n749), .B(datain[3]), .Y(n741) );
  nor4_1 U1012 ( .A(n984), .B(datain[0]), .C(datain[6]), .D(op[1]), .Y(n901)
         );
  nand2_1 U1013 ( .A(n622), .B(n727), .Y(n984) );
  o32ai_1 U1014 ( .A1(n837), .A2(n578), .A3(n924), .B1(n995), .B2(n996), .Y(
        n992) );
  nand2_1 U1015 ( .A(n890), .B(n745), .Y(n996) );
  nor2_1 U1016 ( .A(n749), .B(n910), .Y(n745) );
  inv_1 U1017 ( .A(datain[3]), .Y(n910) );
  inv_1 U1018 ( .A(datain[4]), .Y(n749) );
  inv_1 U1019 ( .A(n856), .Y(n890) );
  nand3_1 U1020 ( .A(n1029), .B(n1031), .C(n989), .Y(n856) );
  inv_1 U1021 ( .A(n941), .Y(n995) );
  nor3_1 U1022 ( .A(n920), .B(datain[0]), .C(n685), .Y(n941) );
  nand2_1 U1023 ( .A(datain[6]), .B(op[1]), .Y(n685) );
  inv_1 U1024 ( .A(n634), .Y(n920) );
  nor2_1 U1025 ( .A(n622), .B(datain[2]), .Y(n634) );
  inv_1 U1026 ( .A(op[0]), .Y(n622) );
  inv_1 U1027 ( .A(n733), .Y(n924) );
  nor3_1 U1028 ( .A(datain[0]), .B(datain[6]), .C(n881), .Y(n733) );
  inv_1 U1029 ( .A(op[1]), .Y(n881) );
  nand2_1 U1030 ( .A(n734), .B(n605), .Y(n578) );
  nor2_1 U1031 ( .A(n727), .B(op[0]), .Y(n605) );
  inv_1 U1032 ( .A(datain[2]), .Y(n727) );
  nor2_1 U1033 ( .A(datain[4]), .B(datain[3]), .Y(n734) );
  nand2_1 U1034 ( .A(n989), .B(n979), .Y(n837) );
  nor2_1 U1035 ( .A(n1029), .B(n1031), .Y(n979) );
  and2_0 U1036 ( .A(n1030), .B(n994), .X(n989) );
  nand2_1 U1037 ( .A(n651), .B(n784), .Y(n994) );
  nor2_1 U1038 ( .A(n1028), .B(n1017), .Y(n784) );
  nor2_1 U1039 ( .A(n1032), .B(n1033), .Y(n651) );
  nor3_1 U1040 ( .A(n998), .B(n997), .C(n1000), .Y(n843) );
endmodule

